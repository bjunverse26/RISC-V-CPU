    rom[0]  = 32'h00500093;
    rom[1]  = 32'h00700113;
    rom[2]  = 32'h002081B3;
    rom[3]  = 32'h00302023;
    rom[4]  = 32'h00002203;
    rom[5]  = 32'h04321463;
    rom[6]  = 32'h123452B7;
    rom[7]  = 32'h00000317;
    rom[8]  = 32'h008003EF;
    rom[9]  = 32'h06300413;
    rom[10] = 32'h02A00413;
    rom[11] = 32'h03400493;
    rom[12] = 32'h00448067;
    rom[13] = 32'h04D00513;
    rom[14] = 32'h00801223;
    rom[15] = 32'h00405583;
    rom[16] = 32'h00100323;
    rom[17] = 32'h00604603;
    rom[18] = 32'h0020C463;
    rom[19] = 32'h00100693;
    rom[20] = 32'h00200693;
    rom[21] = 32'h00D02423;
    rom[22] = 32'h0000006F;
    rom[23] = 32'h07F00693;
    rom[24] = 32'h00D02423;
    rom[25] = 32'h0000006F;
